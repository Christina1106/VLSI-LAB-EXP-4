//MOD -10 COUNTER 
module counter(
input clk,rst, enable,
output reg [3:0]counter_output 
);
always@ (posedge clk)
begin
if(rst | counter_output==4'b1001)
counter_output <= 4'b0000;
else if(enable)
counter_output <= counter_output + 1;
else
counter_output <= 0;
end
endmodule
